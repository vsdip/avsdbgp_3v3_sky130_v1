magic
tech sky130A
magscale 1 2
timestamp 1616724825
<< nwell >>
rect -600 19200 7000 20000
rect -562 17388 -256 19200
rect 1536 18258 5860 19200
rect 1786 18204 5860 18258
rect 1536 15050 5860 18204
<< mvpsubdiff >>
rect -500 4400 6900 4580
rect -500 4200 -440 4400
rect -240 4200 160 4400
rect 360 4200 760 4400
rect 960 4200 1360 4400
rect 1560 4200 1960 4400
rect 2160 4200 2560 4400
rect 2760 4200 3160 4400
rect 3360 4200 3760 4400
rect 3960 4200 4360 4400
rect 4560 4200 4960 4400
rect 5160 4200 5560 4400
rect 5760 4200 6160 4400
rect 6360 4200 6900 4400
rect -500 4020 6900 4200
<< mvnsubdiff >>
rect -500 19700 6900 19880
rect -500 19500 -440 19700
rect -240 19500 160 19700
rect 360 19500 760 19700
rect 960 19500 1360 19700
rect 1560 19500 1960 19700
rect 2160 19500 2560 19700
rect 2760 19500 3160 19700
rect 3360 19500 3760 19700
rect 3960 19500 4360 19700
rect 4560 19500 4960 19700
rect 5160 19500 5560 19700
rect 5760 19500 6160 19700
rect 6360 19500 6900 19700
rect -500 19320 6900 19500
<< mvpsubdiffcont >>
rect -440 4200 -240 4400
rect 160 4200 360 4400
rect 760 4200 960 4400
rect 1360 4200 1560 4400
rect 1960 4200 2160 4400
rect 2560 4200 2760 4400
rect 3160 4200 3360 4400
rect 3760 4200 3960 4400
rect 4360 4200 4560 4400
rect 4960 4200 5160 4400
rect 5560 4200 5760 4400
rect 6160 4200 6360 4400
<< mvnsubdiffcont >>
rect -440 19500 -240 19700
rect 160 19500 360 19700
rect 760 19500 960 19700
rect 1360 19500 1560 19700
rect 1960 19500 2160 19700
rect 2560 19500 2760 19700
rect 3160 19500 3360 19700
rect 3760 19500 3960 19700
rect 4360 19500 4560 19700
rect 4960 19500 5160 19700
rect 5560 19500 5760 19700
rect 6160 19500 6360 19700
<< poly >>
rect 2672 18604 3198 19170
rect 2672 18570 2904 18604
rect 2954 18570 3198 18604
rect 2672 18230 3198 18570
rect 2672 18180 3146 18230
rect 3180 18180 3198 18230
rect 2672 18170 3198 18180
rect 4198 18170 4724 19170
rect 2672 14274 3198 14840
rect 2672 14240 2896 14274
rect 2946 14240 3198 14274
rect 2672 13840 3198 14240
rect 2672 9540 3198 10540
rect 4198 9540 4724 10540
<< polycont >>
rect 2904 18570 2954 18604
rect 3146 18180 3180 18230
rect 1102 15068 1170 15102
rect 2896 14240 2946 14274
rect 1692 13954 1742 13988
rect 528 13678 728 13712
rect -310 5302 -276 5352
<< xpolycontact >>
rect 6360 15574 6430 16006
rect 6042 9222 6112 9654
rect 6042 7040 6112 7472
rect 6360 7040 6430 7472
rect 6678 15574 6748 16006
rect 6678 7040 6748 7472
<< xpolyres >>
rect 6042 7472 6112 9222
rect 6360 7472 6430 15574
rect 6678 7472 6748 15574
<< locali >>
rect -600 19700 7000 19880
rect -600 19500 -440 19700
rect -240 19500 160 19700
rect 360 19500 760 19700
rect 960 19500 1360 19700
rect 1560 19500 1960 19700
rect 2160 19500 2560 19700
rect 2760 19500 3160 19700
rect 3360 19500 3760 19700
rect 3960 19500 4360 19700
rect 4560 19500 4960 19700
rect 5160 19500 5560 19700
rect 5760 19500 6160 19700
rect 6360 19500 7000 19700
rect -600 19320 7000 19500
rect -426 17308 -392 19320
rect 984 18570 2544 18604
rect 2594 18570 2610 18604
rect 984 15752 1018 18570
rect 2690 18120 2724 19320
rect 2780 18570 2796 18604
rect 2846 18570 2904 18604
rect 2954 18570 2978 18604
rect 3146 18230 3180 18246
rect 3146 18120 3180 18180
rect 4216 18120 4250 19320
rect 5742 18120 5776 19320
rect 6358 16006 6432 16008
rect 6358 15574 6360 16006
rect 6430 15804 6432 16006
rect 6676 16006 6750 16008
rect 6676 15804 6678 16006
rect 6430 15770 6678 15804
rect 6430 15574 6432 15770
rect 6358 15572 6432 15574
rect 6676 15574 6678 15770
rect 6748 15574 6750 16006
rect 6676 15572 6750 15574
rect 1254 15104 1288 15152
rect -188 15068 1102 15102
rect 1170 15068 1186 15102
rect 1254 15070 1434 15104
rect -310 5352 -276 5368
rect -426 5154 -392 5204
rect -310 5154 -276 5302
rect -188 5154 -154 15068
rect 1400 14574 1434 15070
rect 1620 15096 1654 15120
rect 1620 15040 1654 15046
rect 3146 15096 3180 15120
rect 3146 15040 3180 15046
rect 4672 15096 4706 15120
rect 4672 15040 4706 15046
rect 1400 14512 1434 14524
rect 616 14240 2896 14274
rect 2946 14240 2962 14274
rect 616 13712 650 14240
rect 1620 13954 1692 13988
rect 1742 13954 1758 13988
rect 1400 13910 1434 13918
rect 512 13678 528 13712
rect 728 13678 744 13712
rect -16 5154 18 5222
rect -426 5120 18 5154
rect 1254 5154 1288 5222
rect 1400 5154 1434 13860
rect 1620 13862 1654 13954
rect 1620 13790 1654 13812
rect 3146 13862 3180 13950
rect 3146 13790 3180 13812
rect 2690 10766 2724 10790
rect 2690 10710 2724 10716
rect 4216 10766 4250 10790
rect 4216 10710 4250 10716
rect 3146 9656 6114 9690
rect 2690 9564 2724 9570
rect 2690 9490 2724 9514
rect 3146 9490 3180 9656
rect 6040 9654 6114 9656
rect 4216 9564 4250 9570
rect 4216 9490 4250 9514
rect 4672 9564 4706 9570
rect 4672 9490 4706 9514
rect 6040 9222 6042 9654
rect 6112 9222 6114 9654
rect 6040 9220 6114 9222
rect 6040 7472 6114 7474
rect 1620 7066 1654 7090
rect 1620 7010 1654 7016
rect 5742 7022 5776 7090
rect 5742 6960 5776 6972
rect 6040 7040 6042 7472
rect 6112 7040 6114 7472
rect 6040 6932 6114 7040
rect 6358 7472 6432 7474
rect 6358 7040 6360 7472
rect 6430 7040 6432 7472
rect 6358 7022 6432 7040
rect 6358 6972 6378 7022
rect 6412 6972 6432 7022
rect 6358 6960 6432 6972
rect 6676 7472 6750 7474
rect 6676 7040 6678 7472
rect 6748 7040 6750 7472
rect 6676 7020 6750 7040
rect 6676 6970 6696 7020
rect 6730 6970 6750 7020
rect 6676 6960 6750 6970
rect 6040 6882 6060 6932
rect 6094 6882 6114 6932
rect 6040 6872 6114 6882
rect 1938 6036 2010 6100
rect 2736 6036 2808 6100
rect 3534 6036 3606 6100
rect 4332 6036 4404 6100
rect 5130 6036 5202 6100
rect 1602 5920 5538 5936
rect 1602 5886 5686 5920
rect 1602 5864 5538 5886
rect 1938 5220 2010 5284
rect 2736 5220 2808 5284
rect 3534 5220 3606 5284
rect 4332 5220 4404 5284
rect 5130 5220 5202 5284
rect 1254 5120 1434 5154
rect 1400 4580 1434 5120
rect 5652 4580 5686 5886
rect -600 4400 7000 4580
rect -600 4200 -440 4400
rect -240 4200 160 4400
rect 360 4200 760 4400
rect 960 4200 1360 4400
rect 1560 4200 1960 4400
rect 2160 4200 2560 4400
rect 2760 4200 3160 4400
rect 3360 4200 3760 4400
rect 3960 4200 4360 4400
rect 4560 4200 4960 4400
rect 5160 4200 5560 4400
rect 5760 4200 6160 4400
rect 6360 4200 7000 4400
rect -600 4020 7000 4200
<< viali >>
rect -440 19500 -240 19700
rect 160 19500 360 19700
rect 760 19500 960 19700
rect 1360 19500 1560 19700
rect 1960 19500 2160 19700
rect 2560 19500 2760 19700
rect 3160 19500 3360 19700
rect 3760 19500 3960 19700
rect 4360 19500 4560 19700
rect 4960 19500 5160 19700
rect 5560 19500 5760 19700
rect 6160 19500 6360 19700
rect 2544 18570 2594 18604
rect 2796 18570 2846 18604
rect 1620 15046 1654 15096
rect 3146 15046 3180 15096
rect 4672 15046 4706 15096
rect 1400 14524 1434 14574
rect 1400 13860 1434 13910
rect 1620 13812 1654 13862
rect 3146 13812 3180 13862
rect 2690 10716 2724 10766
rect 4216 10716 4250 10766
rect 2690 9514 2724 9564
rect 4216 9514 4250 9564
rect 4672 9514 4706 9564
rect 1620 7016 1654 7066
rect 5742 6972 5776 7022
rect 6378 6972 6412 7022
rect 6696 6970 6730 7020
rect 6060 6882 6094 6932
rect -440 4200 -240 4400
rect 160 4200 360 4400
rect 760 4200 960 4400
rect 1360 4200 1560 4400
rect 1960 4200 2160 4400
rect 2560 4200 2760 4400
rect 3160 4200 3360 4400
rect 3760 4200 3960 4400
rect 4360 4200 4560 4400
rect 4960 4200 5160 4400
rect 5560 4200 5760 4400
rect 6160 4200 6360 4400
<< metal1 >>
rect -600 19700 7000 19900
rect -600 19500 -440 19700
rect -240 19500 160 19700
rect 360 19500 760 19700
rect 960 19500 1360 19700
rect 1560 19500 1960 19700
rect 2160 19500 2560 19700
rect 2760 19500 3160 19700
rect 3360 19500 3760 19700
rect 3960 19500 4360 19700
rect 4560 19500 4960 19700
rect 5160 19500 5560 19700
rect 5760 19500 6160 19700
rect 6360 19500 7000 19700
rect -600 19300 7000 19500
rect 2500 18604 2858 18618
rect 2500 18570 2544 18604
rect 2594 18570 2796 18604
rect 2846 18570 2858 18604
rect 2500 18558 2858 18570
rect 1606 15096 1666 15110
rect 1606 15046 1620 15096
rect 1654 15046 1666 15096
rect 1388 14574 1448 14588
rect 1388 14524 1400 14574
rect 1434 14524 1448 14574
rect 1388 13910 1448 14524
rect 1388 13860 1400 13910
rect 1434 13860 1448 13910
rect 1388 13846 1448 13860
rect 1606 13862 1666 15046
rect 1606 13812 1620 13862
rect 1654 13812 1666 13862
rect 1606 13800 1666 13812
rect 3132 15096 3192 15110
rect 3132 15046 3146 15096
rect 3180 15046 3192 15096
rect 3132 13862 3192 15046
rect 3132 13812 3146 13862
rect 3180 13812 3192 13862
rect 3132 13800 3192 13812
rect 4658 15096 4718 15110
rect 4658 15046 4672 15096
rect 4706 15046 4718 15096
rect 2678 10766 2738 10780
rect 2678 10716 2690 10766
rect 2724 10716 2738 10766
rect 2678 9564 2738 10716
rect 2678 9514 2690 9564
rect 2724 9514 2738 9564
rect 2678 9500 2738 9514
rect 4204 10766 4264 10780
rect 4204 10716 4216 10766
rect 4250 10716 4264 10766
rect 4204 9564 4264 10716
rect 4204 9514 4216 9564
rect 4250 9514 4264 9564
rect 4204 9500 4264 9514
rect 4658 9564 4718 15046
rect 4658 9514 4672 9564
rect 4706 9514 4718 9564
rect 4658 9500 4718 9514
rect 1606 7066 1666 7080
rect 1606 7016 1620 7066
rect 1654 7016 1666 7066
rect 1606 6886 1666 7016
rect 5730 7022 6424 7028
rect 5730 6972 5742 7022
rect 5776 6972 6378 7022
rect 6412 6972 6424 7022
rect 5730 6966 6424 6972
rect 6682 7020 6742 7032
rect 6682 6970 6696 7020
rect 6730 6970 6742 7020
rect 3540 6932 6114 6938
rect 1606 6826 2004 6886
rect 1944 6390 2004 6826
rect 3540 6882 6060 6932
rect 6094 6882 6114 6932
rect 3540 6876 6114 6882
rect 3540 6790 3600 6876
rect 2316 6730 5196 6790
rect 2316 5522 2376 6730
rect 2742 6390 2802 6730
rect 3114 5522 3174 6730
rect 3540 6390 3600 6730
rect 3912 5522 3972 6730
rect 4338 6390 4398 6730
rect 4710 5522 4770 6730
rect 5136 6390 5196 6730
rect 6682 5522 6742 6970
rect 2056 5462 2376 5522
rect 2854 5462 3174 5522
rect 3652 5462 3972 5522
rect 4450 5462 4770 5522
rect 5248 5462 6742 5522
rect -600 4400 7000 4800
rect -600 4200 -440 4400
rect -240 4200 160 4400
rect 360 4200 760 4400
rect 960 4200 1360 4400
rect 1560 4200 1960 4400
rect 2160 4200 2560 4400
rect 2760 4200 3160 4400
rect 3360 4200 3760 4400
rect 3960 4200 4360 4400
rect 4560 4200 4960 4400
rect 5160 4200 5560 4400
rect 5760 4200 6160 4400
rect 6360 4200 7000 4400
rect -600 3800 7000 4200
use sc_pmos  sc_pmos_0
timestamp 1616540248
transform 1 0 -960 0 1 2192
box 400 2928 700 15200
use sc_nmos_426  sc_nmos_426_0
timestamp 1616700505
transform 1 0 -414 0 1 4020
box 380 1100 1720 9704
use sc_nmos_31  sc_nmos_31_0
timestamp 1616174596
transform 1 0 586 0 1 13950
box 380 1100 720 1904
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1615375237
transform 1 0 1576 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1615375237
transform 1 0 1576 0 1 5094
box 26 26 770 795
use cm_nmos  cm_nmos_1
timestamp 1616067151
transform 1 0 1672 0 1 10740
box -70 0 1070 4100
use en_nmos  en_nmos_0
timestamp 1616065709
transform 1 0 1672 0 1 7040
box -70 0 1070 3500
use cm_pmos  cm_pmos_0
timestamp 1616078161
transform 1 0 1672 0 1 15070
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1615375237
transform 1 0 2374 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1615375237
transform 1 0 2374 0 1 5094
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1615375237
transform 1 0 3172 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1615375237
transform 1 0 3172 0 1 5094
box 26 26 770 795
use en_nmos  en_nmos_1
timestamp 1616065709
transform 1 0 3198 0 1 7040
box -70 0 1070 3500
use cm_nmos  cm_nmos_0
timestamp 1616067151
transform 1 0 3198 0 1 10740
box -70 0 1070 4100
use cm_pmos  cm_pmos_1
timestamp 1616078161
transform 1 0 3198 0 1 15070
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1615375237
transform 1 0 3970 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1615375237
transform 1 0 3970 0 1 5094
box 26 26 770 795
use en_nmos  en_nmos_2
timestamp 1616065709
transform 1 0 4724 0 1 7040
box -70 0 1070 3500
use cm_pmos  cm_pmos_2
timestamp 1616078161
transform 1 0 4724 0 1 15070
box -136 -20 1136 4100
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8
timestamp 1615375237
transform 1 0 4768 0 1 5910
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_9
timestamp 1615375237
transform 1 0 4768 0 1 5094
box 26 26 770 795
<< labels >>
flabel poly s 2754 10146 3176 10506 0 FreeSans 1600 0 0 0 en
flabel locali s 6422 6962 6432 6966 0 FreeSans 400 0 0 0 Vbgp
flabel metal1 s 5896 6886 5954 6902 0 FreeSans 400 0 0 0 A
flabel locali s 5900 9662 5958 9678 0 FreeSans 400 0 0 0 B
flabel metal1 s 4216 10642 4274 10658 0 FreeSans 400 0 0 0 C
flabel metal1 s 3168 14956 3226 14972 0 FreeSans 400 0 0 0 D
flabel metal1 s 4694 14940 4708 14960 0 FreeSans 400 0 0 0 E
flabel metal1 s 1646 6976 1660 6996 0 FreeSans 400 0 0 0 F
flabel metal1 s 2704 10660 2718 10680 0 FreeSans 400 0 0 0 G
flabel locali s 6534 15786 6548 15806 0 FreeSans 400 0 0 0 H
flabel metal1 s 6702 6792 6716 6812 0 FreeSans 400 0 0 0 J
flabel locali s -184 5124 -176 5130 0 FreeSans 800 0 0 0 I
flabel locali s 712 14256 722 14266 0 FreeSans 800 0 0 0 VbiasN
flabel locali s 1028 18590 1038 18598 0 FreeSans 800 0 0 0 VbiasP
flabel locali s -346 4056 -332 4072 0 FreeSans 800 0 0 0 GND
flabel locali s -362 19764 -348 19780 0 FreeSans 800 0 0 0 VDD
<< end >>
