magic
tech sky130A
timestamp 1616540248
<< nwell >>
rect 200 1464 350 7600
<< mvpmos >>
rect 250 1532 300 7532
<< mvpdiff >>
rect 250 7558 300 7567
rect 250 7541 258 7558
rect 292 7541 300 7558
rect 250 7532 300 7541
rect 250 1523 300 1532
rect 250 1506 258 1523
rect 292 1506 300 1523
rect 250 1497 300 1506
<< mvpdiffc >>
rect 258 7541 292 7558
rect 258 1506 292 1523
<< poly >>
rect 200 1532 250 7532
rect 300 1532 350 7532
<< locali >>
rect 250 7541 258 7558
rect 292 7541 300 7558
rect 250 1506 258 1523
rect 292 1506 300 1523
<< end >>
