magic
tech sky130A
timestamp 1616067151
<< mvnmos >>
rect 0 25 500 1525
<< mvndiff >>
rect -35 1485 0 1525
rect -35 1385 -26 1485
rect -9 1385 0 1485
rect -35 1365 0 1385
rect -35 1265 -26 1365
rect -9 1265 0 1365
rect -35 1245 0 1265
rect -35 1145 -26 1245
rect -9 1145 0 1245
rect -35 1125 0 1145
rect -35 1025 -26 1125
rect -9 1025 0 1125
rect -35 1005 0 1025
rect -35 905 -26 1005
rect -9 905 0 1005
rect -35 885 0 905
rect -35 785 -26 885
rect -9 785 0 885
rect -35 765 0 785
rect -35 665 -26 765
rect -9 665 0 765
rect -35 645 0 665
rect -35 545 -26 645
rect -9 545 0 645
rect -35 525 0 545
rect -35 425 -26 525
rect -9 425 0 525
rect -35 405 0 425
rect -35 305 -26 405
rect -9 305 0 405
rect -35 285 0 305
rect -35 185 -26 285
rect -9 185 0 285
rect -35 165 0 185
rect -35 65 -26 165
rect -9 65 0 165
rect -35 25 0 65
rect 500 1485 535 1525
rect 500 1385 509 1485
rect 526 1385 535 1485
rect 500 1365 535 1385
rect 500 1265 509 1365
rect 526 1265 535 1365
rect 500 1245 535 1265
rect 500 1145 509 1245
rect 526 1145 535 1245
rect 500 1125 535 1145
rect 500 1025 509 1125
rect 526 1025 535 1125
rect 500 1005 535 1025
rect 500 905 509 1005
rect 526 905 535 1005
rect 500 885 535 905
rect 500 785 509 885
rect 526 785 535 885
rect 500 765 535 785
rect 500 665 509 765
rect 526 665 535 765
rect 500 645 535 665
rect 500 545 509 645
rect 526 545 535 645
rect 500 525 535 545
rect 500 425 509 525
rect 526 425 535 525
rect 500 405 535 425
rect 500 305 509 405
rect 526 305 535 405
rect 500 285 535 305
rect 500 185 509 285
rect 526 185 535 285
rect 500 165 535 185
rect 500 65 509 165
rect 526 65 535 165
rect 500 25 535 65
<< mvndiffc >>
rect -26 1385 -9 1485
rect -26 1265 -9 1365
rect -26 1145 -9 1245
rect -26 1025 -9 1125
rect -26 905 -9 1005
rect -26 785 -9 885
rect -26 665 -9 765
rect -26 545 -9 645
rect -26 425 -9 525
rect -26 305 -9 405
rect -26 185 -9 285
rect -26 65 -9 165
rect 509 1385 526 1485
rect 509 1265 526 1365
rect 509 1145 526 1245
rect 509 1025 526 1125
rect 509 905 526 1005
rect 509 785 526 885
rect 509 665 526 765
rect 509 545 526 645
rect 509 425 526 525
rect 509 305 526 405
rect 509 185 526 285
rect 509 65 526 165
<< poly >>
rect 0 1525 500 2050
rect 0 0 500 25
<< locali >>
rect -26 1485 -9 1525
rect -26 1365 -9 1385
rect -26 1245 -9 1265
rect -26 1125 -9 1145
rect -26 1005 -9 1025
rect -26 885 -9 905
rect -26 765 -9 785
rect -26 645 -9 665
rect -26 525 -9 545
rect -26 405 -9 425
rect -26 285 -9 305
rect -26 165 -9 185
rect -26 25 -9 65
rect 509 1485 526 1525
rect 509 1365 526 1385
rect 509 1245 526 1265
rect 509 1125 526 1145
rect 509 1005 526 1025
rect 509 885 526 905
rect 509 765 526 785
rect 509 645 526 665
rect 509 525 526 545
rect 509 405 526 425
rect 509 285 526 305
rect 509 165 526 185
rect 509 25 526 65
<< end >>
