magic
tech sky130A
timestamp 1616065709
<< mvnmos >>
rect 0 25 500 1225
<< mvndiff >>
rect -35 1215 0 1225
rect -35 1115 -26 1215
rect -9 1115 0 1215
rect -35 1095 0 1115
rect -35 995 -26 1095
rect -9 995 0 1095
rect -35 975 0 995
rect -35 875 -26 975
rect -9 875 0 975
rect -35 855 0 875
rect -35 755 -26 855
rect -9 755 0 855
rect -35 735 0 755
rect -35 635 -26 735
rect -9 635 0 735
rect -35 615 0 635
rect -35 515 -26 615
rect -9 515 0 615
rect -35 495 0 515
rect -35 395 -26 495
rect -9 395 0 495
rect -35 375 0 395
rect -35 275 -26 375
rect -9 275 0 375
rect -35 255 0 275
rect -35 155 -26 255
rect -9 155 0 255
rect -35 135 0 155
rect -35 35 -26 135
rect -9 35 0 135
rect -35 25 0 35
rect 500 1215 535 1225
rect 500 1115 509 1215
rect 526 1115 535 1215
rect 500 1095 535 1115
rect 500 995 509 1095
rect 526 995 535 1095
rect 500 975 535 995
rect 500 875 509 975
rect 526 875 535 975
rect 500 855 535 875
rect 500 755 509 855
rect 526 755 535 855
rect 500 735 535 755
rect 500 635 509 735
rect 526 635 535 735
rect 500 615 535 635
rect 500 515 509 615
rect 526 515 535 615
rect 500 495 535 515
rect 500 395 509 495
rect 526 395 535 495
rect 500 375 535 395
rect 500 275 509 375
rect 526 275 535 375
rect 500 255 535 275
rect 500 155 509 255
rect 526 155 535 255
rect 500 135 535 155
rect 500 35 509 135
rect 526 35 535 135
rect 500 25 535 35
<< mvndiffc >>
rect -26 1115 -9 1215
rect -26 995 -9 1095
rect -26 875 -9 975
rect -26 755 -9 855
rect -26 635 -9 735
rect -26 515 -9 615
rect -26 395 -9 495
rect -26 275 -9 375
rect -26 155 -9 255
rect -26 35 -9 135
rect 509 1115 526 1215
rect 509 995 526 1095
rect 509 875 526 975
rect 509 755 526 855
rect 509 635 526 735
rect 509 515 526 615
rect 509 395 526 495
rect 509 275 526 375
rect 509 155 526 255
rect 509 35 526 135
<< poly >>
rect 0 1225 500 1750
rect 0 0 500 25
<< locali >>
rect -26 1215 -9 1225
rect -26 1095 -9 1115
rect -26 975 -9 995
rect -26 855 -9 875
rect -26 735 -9 755
rect -26 615 -9 635
rect -26 495 -9 515
rect -26 375 -9 395
rect -26 255 -9 275
rect -26 135 -9 155
rect -26 25 -9 35
rect 509 1215 526 1225
rect 509 1095 526 1115
rect 509 975 526 995
rect 509 855 526 875
rect 509 735 526 755
rect 509 615 526 635
rect 509 495 526 515
rect 509 375 526 395
rect 509 255 526 275
rect 509 135 526 155
rect 509 25 526 35
<< end >>
