magic
tech sky130A
timestamp 1616174596
<< mvnmos >>
rect 225 601 325 901
<< mvndiff >>
rect 190 892 225 901
rect 190 801 199 892
rect 216 801 225 892
rect 190 701 225 801
rect 190 610 199 701
rect 216 610 225 701
rect 190 601 225 610
rect 325 892 360 901
rect 325 801 334 892
rect 351 801 360 892
rect 325 701 360 801
rect 325 610 334 701
rect 351 610 360 701
rect 325 601 360 610
<< mvndiffc >>
rect 199 801 216 892
rect 199 610 216 701
rect 334 801 351 892
rect 334 610 351 701
<< poly >>
rect 225 901 325 952
rect 225 550 325 601
<< locali >>
rect 199 892 216 901
rect 199 701 216 801
rect 199 601 216 610
rect 334 892 351 901
rect 334 701 351 801
rect 334 601 351 610
<< end >>
