**.subckt avsdbgp_3V3
XM1 VbiasN VbiasN net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 VbiasP VbiasN net4 GND sky130_fd_pr__nfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 VbiasN VbiasP VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XQ1 GND GND Vleft_branch GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ2 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XM5 net2 VbiasP VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XQ3 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ4 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ5 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ6 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ7 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ8 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XQ9 GND GND net1 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
R1 Vright_branch net1 50k m=1
R2 Vbgp net6 463k m=1
XQ10 GND GND net6 GND sky130_fd_pr__pnp_05v5_W3p40L3p40
XM4 VbiasP VbiasP VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=15 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7 net5 VbiasN GND GND sky130_fd_pr__nfet_g5v0d10v5 L=6 W=42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 VbiasP net5 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
RLoad Vbgp GND 100Meg m=1
XM9 net3 en Vleft_branch GND sky130_fd_pr__nfet_g5v0d10v5 L=5 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM10 net4 en Vright_branch GND sky130_fd_pr__nfet_g5v0d10v5 L=5 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM11 net2 en Vbgp GND sky130_fd_pr__nfet_g5v0d10v5 L=5 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 net5 net5 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=60 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
**** begin user architecture code


.lib ../../lib/models/sky130_tt_bgr.lib.spice tt
.options savecurrents

*** plot vbgp with variation in supply voltage
*Vdd VDD GND 3.3
*V_en en GND 3.3
*.dc Vdd 2 4 0.1
*.control
*run
*print Vbgp
*plot V(Vbgp)
*.endc

*** plot vbgp with variation in temperature @3.3V
*Vdd VDD GND 3.3
*V_en en GND 3.3
*.dc temp -40 140 1
*.control
*run
*print V(Vbgp)
*plot V(Vbgp)
*.endc

*** plot voltage coefficient
*Vdd VDD GND 3.3
*V_en en GND 3.3
*.dc Vdd 2 4 0.1
*.control
*run
*plot deriv(V(Vbgp))
*.endc

*** plot temperature coefficient
*Vdd VDD GND 3.3
*V_en en GND 3.3
*.dc temp -40 140 1
*.control
*run
*plot deriv(V(Vbgp))/1.202344
*.endc

*** check start up circuit
V_en en GND 3.3
Vdd VDD GND PULSE(0 3.3 50us 200us 200us 600us 2000us 0)
.tran 1us 800us
.control
run
plot V(Vdd) V(Vbgp)
.endc

*** enable pin
*Vdd VDD GND 3.3
*V_en en GND PULSE(0 3.3 0 2000us 2000us 6000us 20000us 0)
*.tran 1u 20000us
*.control
*run
*plot V(en)
*plot -I(VDD)
*.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.GLOBAL en
** flattened .save nodes
.end
