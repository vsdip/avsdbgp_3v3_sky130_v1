magic
tech sky130A
timestamp 1616700505
<< mvnmos >>
rect 225 601 825 4801
<< mvndiff >>
rect 190 4790 225 4801
rect 190 4690 199 4790
rect 216 4690 225 4790
rect 190 4670 225 4690
rect 190 4570 199 4670
rect 216 4570 225 4670
rect 190 4550 225 4570
rect 190 4450 199 4550
rect 216 4450 225 4550
rect 190 4430 225 4450
rect 190 4330 199 4430
rect 216 4330 225 4430
rect 190 4310 225 4330
rect 190 4210 199 4310
rect 216 4210 225 4310
rect 190 4190 225 4210
rect 190 4090 199 4190
rect 216 4090 225 4190
rect 190 4070 225 4090
rect 190 3970 199 4070
rect 216 3970 225 4070
rect 190 3950 225 3970
rect 190 3850 199 3950
rect 216 3850 225 3950
rect 190 3830 225 3850
rect 190 3730 199 3830
rect 216 3730 225 3830
rect 190 3710 225 3730
rect 190 3610 199 3710
rect 216 3610 225 3710
rect 190 3590 225 3610
rect 190 3490 199 3590
rect 216 3490 225 3590
rect 190 3470 225 3490
rect 190 3370 199 3470
rect 216 3370 225 3470
rect 190 3350 225 3370
rect 190 3250 199 3350
rect 216 3250 225 3350
rect 190 3230 225 3250
rect 190 3130 199 3230
rect 216 3130 225 3230
rect 190 3110 225 3130
rect 190 3010 199 3110
rect 216 3010 225 3110
rect 190 2990 225 3010
rect 190 2890 199 2990
rect 216 2890 225 2990
rect 190 2870 225 2890
rect 190 2770 199 2870
rect 216 2770 225 2870
rect 190 2750 225 2770
rect 190 2650 199 2750
rect 216 2650 225 2750
rect 190 2630 225 2650
rect 190 2530 199 2630
rect 216 2530 225 2630
rect 190 2510 225 2530
rect 190 2410 199 2510
rect 216 2410 225 2510
rect 190 2390 225 2410
rect 190 2290 199 2390
rect 216 2290 225 2390
rect 190 2270 225 2290
rect 190 2170 199 2270
rect 216 2170 225 2270
rect 190 2150 225 2170
rect 190 2050 199 2150
rect 216 2050 225 2150
rect 190 2030 225 2050
rect 190 1930 199 2030
rect 216 1930 225 2030
rect 190 1910 225 1930
rect 190 1810 199 1910
rect 216 1810 225 1910
rect 190 1790 225 1810
rect 190 1690 199 1790
rect 216 1690 225 1790
rect 190 1670 225 1690
rect 190 1570 199 1670
rect 216 1570 225 1670
rect 190 1550 225 1570
rect 190 1450 199 1550
rect 216 1450 225 1550
rect 190 1430 225 1450
rect 190 1330 199 1430
rect 216 1330 225 1430
rect 190 1310 225 1330
rect 190 1210 199 1310
rect 216 1210 225 1310
rect 190 1190 225 1210
rect 190 1090 199 1190
rect 216 1090 225 1190
rect 190 1070 225 1090
rect 190 970 199 1070
rect 216 970 225 1070
rect 190 950 225 970
rect 190 850 199 950
rect 216 850 225 950
rect 190 830 225 850
rect 190 730 199 830
rect 216 730 225 830
rect 190 710 225 730
rect 190 610 199 710
rect 216 610 225 710
rect 190 601 225 610
rect 825 4790 860 4801
rect 825 4690 834 4790
rect 851 4690 860 4790
rect 825 4670 860 4690
rect 825 4570 834 4670
rect 851 4570 860 4670
rect 825 4550 860 4570
rect 825 4450 834 4550
rect 851 4450 860 4550
rect 825 4430 860 4450
rect 825 4330 834 4430
rect 851 4330 860 4430
rect 825 4310 860 4330
rect 825 4210 834 4310
rect 851 4210 860 4310
rect 825 4190 860 4210
rect 825 4090 834 4190
rect 851 4090 860 4190
rect 825 4070 860 4090
rect 825 3970 834 4070
rect 851 3970 860 4070
rect 825 3950 860 3970
rect 825 3850 834 3950
rect 851 3850 860 3950
rect 825 3830 860 3850
rect 825 3730 834 3830
rect 851 3730 860 3830
rect 825 3710 860 3730
rect 825 3610 834 3710
rect 851 3610 860 3710
rect 825 3590 860 3610
rect 825 3490 834 3590
rect 851 3490 860 3590
rect 825 3470 860 3490
rect 825 3370 834 3470
rect 851 3370 860 3470
rect 825 3350 860 3370
rect 825 3250 834 3350
rect 851 3250 860 3350
rect 825 3230 860 3250
rect 825 3130 834 3230
rect 851 3130 860 3230
rect 825 3110 860 3130
rect 825 3010 834 3110
rect 851 3010 860 3110
rect 825 2990 860 3010
rect 825 2890 834 2990
rect 851 2890 860 2990
rect 825 2870 860 2890
rect 825 2770 834 2870
rect 851 2770 860 2870
rect 825 2750 860 2770
rect 825 2650 834 2750
rect 851 2650 860 2750
rect 825 2630 860 2650
rect 825 2530 834 2630
rect 851 2530 860 2630
rect 825 2510 860 2530
rect 825 2410 834 2510
rect 851 2410 860 2510
rect 825 2390 860 2410
rect 825 2290 834 2390
rect 851 2290 860 2390
rect 825 2270 860 2290
rect 825 2170 834 2270
rect 851 2170 860 2270
rect 825 2150 860 2170
rect 825 2050 834 2150
rect 851 2050 860 2150
rect 825 2030 860 2050
rect 825 1930 834 2030
rect 851 1930 860 2030
rect 825 1910 860 1930
rect 825 1810 834 1910
rect 851 1810 860 1910
rect 825 1790 860 1810
rect 825 1690 834 1790
rect 851 1690 860 1790
rect 825 1670 860 1690
rect 825 1570 834 1670
rect 851 1570 860 1670
rect 825 1550 860 1570
rect 825 1450 834 1550
rect 851 1450 860 1550
rect 825 1430 860 1450
rect 825 1330 834 1430
rect 851 1330 860 1430
rect 825 1310 860 1330
rect 825 1210 834 1310
rect 851 1210 860 1310
rect 825 1190 860 1210
rect 825 1090 834 1190
rect 851 1090 860 1190
rect 825 1070 860 1090
rect 825 970 834 1070
rect 851 970 860 1070
rect 825 950 860 970
rect 825 850 834 950
rect 851 850 860 950
rect 825 830 860 850
rect 825 730 834 830
rect 851 730 860 830
rect 825 710 860 730
rect 825 610 834 710
rect 851 610 860 710
rect 825 601 860 610
<< mvndiffc >>
rect 199 4690 216 4790
rect 199 4570 216 4670
rect 199 4450 216 4550
rect 199 4330 216 4430
rect 199 4210 216 4310
rect 199 4090 216 4190
rect 199 3970 216 4070
rect 199 3850 216 3950
rect 199 3730 216 3830
rect 199 3610 216 3710
rect 199 3490 216 3590
rect 199 3370 216 3470
rect 199 3250 216 3350
rect 199 3130 216 3230
rect 199 3010 216 3110
rect 199 2890 216 2990
rect 199 2770 216 2870
rect 199 2650 216 2750
rect 199 2530 216 2630
rect 199 2410 216 2510
rect 199 2290 216 2390
rect 199 2170 216 2270
rect 199 2050 216 2150
rect 199 1930 216 2030
rect 199 1810 216 1910
rect 199 1690 216 1790
rect 199 1570 216 1670
rect 199 1450 216 1550
rect 199 1330 216 1430
rect 199 1210 216 1310
rect 199 1090 216 1190
rect 199 970 216 1070
rect 199 850 216 950
rect 199 730 216 830
rect 199 610 216 710
rect 834 4690 851 4790
rect 834 4570 851 4670
rect 834 4450 851 4550
rect 834 4330 851 4430
rect 834 4210 851 4310
rect 834 4090 851 4190
rect 834 3970 851 4070
rect 834 3850 851 3950
rect 834 3730 851 3830
rect 834 3610 851 3710
rect 834 3490 851 3590
rect 834 3370 851 3470
rect 834 3250 851 3350
rect 834 3130 851 3230
rect 834 3010 851 3110
rect 834 2890 851 2990
rect 834 2770 851 2870
rect 834 2650 851 2750
rect 834 2530 851 2630
rect 834 2410 851 2510
rect 834 2290 851 2390
rect 834 2170 851 2270
rect 834 2050 851 2150
rect 834 1930 851 2030
rect 834 1810 851 1910
rect 834 1690 851 1790
rect 834 1570 851 1670
rect 834 1450 851 1550
rect 834 1330 851 1430
rect 834 1210 851 1310
rect 834 1090 851 1190
rect 834 970 851 1070
rect 834 850 851 950
rect 834 730 851 830
rect 834 610 851 710
<< poly >>
rect 225 4801 825 4852
rect 225 550 825 601
<< locali >>
rect 199 4790 216 4801
rect 199 4670 216 4690
rect 199 4550 216 4570
rect 199 4430 216 4450
rect 199 4310 216 4330
rect 199 4190 216 4210
rect 199 4070 216 4090
rect 199 3950 216 3970
rect 199 3830 216 3850
rect 199 3710 216 3730
rect 199 3590 216 3610
rect 199 3470 216 3490
rect 199 3350 216 3370
rect 199 3230 216 3250
rect 199 3110 216 3130
rect 199 2990 216 3010
rect 199 2870 216 2890
rect 199 2750 216 2770
rect 199 2630 216 2650
rect 199 2510 216 2530
rect 199 2390 216 2410
rect 199 2270 216 2290
rect 199 2150 216 2170
rect 199 2030 216 2050
rect 199 1910 216 1930
rect 199 1790 216 1810
rect 199 1670 216 1690
rect 199 1550 216 1570
rect 199 1430 216 1450
rect 199 1310 216 1330
rect 199 1190 216 1210
rect 199 1070 216 1090
rect 199 950 216 970
rect 199 830 216 850
rect 199 710 216 730
rect 199 601 216 610
rect 834 4790 851 4801
rect 834 4670 851 4690
rect 834 4550 851 4570
rect 834 4430 851 4450
rect 834 4310 851 4330
rect 834 4190 851 4210
rect 834 4070 851 4090
rect 834 3950 851 3970
rect 834 3830 851 3850
rect 834 3710 851 3730
rect 834 3590 851 3610
rect 834 3470 851 3490
rect 834 3350 851 3370
rect 834 3230 851 3250
rect 834 3110 851 3130
rect 834 2990 851 3010
rect 834 2870 851 2890
rect 834 2750 851 2770
rect 834 2630 851 2650
rect 834 2510 851 2530
rect 834 2390 851 2410
rect 834 2270 851 2290
rect 834 2150 851 2170
rect 834 2030 851 2050
rect 834 1910 851 1930
rect 834 1790 851 1810
rect 834 1670 851 1690
rect 834 1550 851 1570
rect 834 1430 851 1450
rect 834 1310 851 1330
rect 834 1190 851 1210
rect 834 1070 851 1090
rect 834 950 851 970
rect 834 830 851 850
rect 834 710 851 730
rect 834 601 851 610
<< end >>
